module flash_control (
	input logic clk,
	input logic rst,
	
	input logic save,
	input logic read,

	output save_req_a,
	output save_req_v,
	input  save_req_d
);

endmodule
