module res_divider (
    input real v_in,
    output real v_out_10
    output real v_out_100
    output real v_out_1000
    output real v_out_10000
);

endmodule