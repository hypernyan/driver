parameter int ADDR_FREQ     = 0;
parameter int ADDR_DUTY     = 1;
parameter int ADDR_PHASE    = 2;
parameter int ADDR_OCD      = 3;
parameter int ADDR_DEADTIME = 4;
parameter int ADDR_CURRENT  = 5;
parameter int ADDR_MOD_FREQ  = 6;
parameter int ADDR_STOP     = ADDR_CURRENT;